module booth (
    input logic clk,
    input logic rst,
    input logic [31:0] multiplicand,
    input logic [31:0] multiplier,
    output logic [63:0] product,
    output logic ready,
);

    
endmodule