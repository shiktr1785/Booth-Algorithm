module mult11s8s (
    clk,        //Declare the design module
    n1,
    n2,
    result
);

input clk;      //Declare the input and output ports
input [10:0] n1;
input [7:0] n2;
output [18:0] result;

//Declare Combination Circuit
wire n1orn2z;
wire [10:0] p1;
wire [10:0] p2;
wire [10:0] p3;
wire [10:0] p4;
wire [10:0] p5;
wire [10:0] p6;
wire [10:0] p7;
wire [10:0] p8;

wire [6:0] s11a;
wire [6:0] s12a;


endmodule